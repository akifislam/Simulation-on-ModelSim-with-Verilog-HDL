module ThreeBitSynchronousUpCounter(Q)
